/icd/ssv_pe_t3/general_timing/aayushis/PARADIME_RAK/libs/lef/FreePDK45_lib_v1.0.lef