/icd/ssv_pe_t3/general_timing/aayushis/PARADIME_RAK/libs/MACRO/LEF/pllclk.lef